-------------------------------------------------
--  File:          InstructionMemory.vhd
--
--  Entity:        InstructionMemory
--  Architecture:  idk
--  Author:        Trent Wesley
--  Created:       02/10/22
--  VHDL'93
--  Description:   The following is the entity and
--                 architectural description of 
--                 instruction memory
-------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity InstructionMemory is
    port (
        addr : in std_logic_vector(27 downto 0);
        d_out : out std_logic_vector(31 downto 0));
end entity InstructionMemory;

architecture idk of InstructionMemory is
    type mem is array (0 to 1023) of std_logic_vector(7 downto 0);
    signal mem_array : mem := (
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"34", x"21", x"00", x"04", -- ORI  $1,$1,4
        x"34", x"42", x"00", x"05", -- ORI  $2,$2,5
        x"34", x"E7", x"00", x"02", -- ORI  $7,$7,2 
        x"35", x"08", x"00", x"02", -- ORI  $8,$8,2 
        x"35", x"29", x"F0", x"00", -- ORI  $9,$9,2 
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", 
        x"00", x"41", x"18", x"20", -- ADD  $3,$2,$1
        x"00", x"41", x"20", x"24", -- AND  $4,$2,$1
        x"00", x"41", x"28", x"19", -- MULTU $5,$2,%1 
        x"00", x"22", x"30", x"25", -- OR   $6,$1,$2
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"00", x"E7", x"38", x"00", -- SLL  $7,$7,$7
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"00", x"E8", x"38", x"02", -- SRL  $7,$7,$8
        x"01", x"28", x"48", x"03", -- SRA  $9,$9,$8
        x"00", x"23", x"08", x"22", -- SUB  $1,$1,$3
        x"00", x"C4", x"30", x"26", -- XOR  $6,$6,$4
        x"20", x"63", x"00", x"07", -- ADDI $3,$3,7
        x"30", x"E7", x"FF", x"FD", -- ANDI $7,$7,0xFFFD
        x"38", x"AA", x"12", x"34", -- XORI $10,$5,0x1234
        x"AD", x"64", x"00", x"14", -- SW   $4,20($11)
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"8D", x"6B", x"00", x"14", -- LW   $11,20($11)
        
        --Fibonacci Start
        x"36", x"94", x"03", x"FF", -- ORI  $20,$20,0x3FF
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"36", x"B5", x"00", x"01", -- ORI  $21,$21,1
        x"AE", x"96", x"00", x"00", -- SW  $22,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"AE", x"95", x"00", x"00", -- SW  $21,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        --1
        x"32", x"F7", x"00", x"00", -- ANDI $23,$23,0
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"F5", x"B8", x"25", -- OR   $23,$23,$21
        x"02", x"B6", x"A8", x"20", -- ADD  $21,$21,$22
        x"32", x"D6", x"00", x"00", -- ANDI $22,$22,0 
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"D7", x"B0", x"25", -- OR   $22,$22,$23 
        x"AE", x"95", x"00", x"00", -- SW  $21,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        --2
        x"32", x"F7", x"00", x"00", -- ANDI $23,$23,0
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"F5", x"B8", x"25", -- OR   $23,$23,$21
        x"02", x"B6", x"A8", x"20", -- ADD  $21,$21,$22
        x"32", x"D6", x"00", x"00", -- ANDI $22,$22,0 
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"D7", x"B0", x"25", -- OR   $22,$22,$23
        x"AE", x"95", x"00", x"00", -- SW  $21,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        --3
        x"32", x"F7", x"00", x"00", -- ANDI $23,$23,0
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"F5", x"B8", x"25", -- OR   $23,$23,$21
        x"02", x"B6", x"A8", x"20", -- ADD  $21,$21,$22
        x"32", x"D6", x"00", x"00", -- ANDI $22,$22,0 
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"D7", x"B0", x"25", -- OR   $22,$22,$23 
        x"AE", x"95", x"00", x"00", -- SW  $21,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        --4
        x"32", x"F7", x"00", x"00", -- ANDI $23,$23,0
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"F5", x"B8", x"25", -- OR   $23,$23,$21
        x"02", x"B6", x"A8", x"20", -- ADD  $21,$21,$22
        x"32", x"D6", x"00", x"00", -- ANDI $22,$22,0 
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"D7", x"B0", x"25", -- OR   $22,$22,$23  
        x"AE", x"95", x"00", x"00", -- SW  $21,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        --5
        x"32", x"F7", x"00", x"00", -- ANDI $23,$23,0
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"F5", x"B8", x"25", -- OR   $23,$23,$21
        x"02", x"B6", x"A8", x"20", -- ADD  $21,$21,$22
        x"32", x"D6", x"00", x"00", -- ANDI $22,$22,0 
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"D7", x"B0", x"25", -- OR   $22,$22,$23
        x"AE", x"95", x"00", x"00", -- SW  $21,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        --6 
        x"32", x"F7", x"00", x"00", -- ANDI $23,$23,0
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"F5", x"B8", x"25", -- OR   $23,$23,$21
        x"02", x"B6", x"A8", x"20", -- ADD  $21,$21,$22
        x"32", x"D6", x"00", x"00", -- ANDI $22,$22,0 
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"D7", x"B0", x"25", -- OR   $22,$22,$23
        x"AE", x"95", x"00", x"00", -- SW  $21,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        --7 
        x"32", x"F7", x"00", x"00", -- ANDI $23,$23,0
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"F5", x"B8", x"25", -- OR   $23,$23,$21
        x"02", x"B6", x"A8", x"20", -- ADD  $21,$21,$22
        x"32", x"D6", x"00", x"00", -- ANDI $22,$22,0 
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"D7", x"B0", x"25", -- OR   $22,$22,$23 
        x"AE", x"95", x"00", x"00", -- SW  $21,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        --8 
        x"32", x"F7", x"00", x"00", -- ANDI $23,$23,0
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"F5", x"B8", x"25", -- OR   $23,$23,$21
        x"02", x"B6", x"A8", x"20", -- ADD  $21,$21,$22
        x"32", x"D6", x"00", x"00", -- ANDI $22,$22,0 
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"D7", x"B0", x"25", -- OR   $22,$22,$23 
        x"AE", x"95", x"00", x"00", -- SW  $21,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        --9 
        x"32", x"F7", x"00", x"00", -- ANDI $23,$23,0
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"F5", x"B8", x"25", -- OR   $23,$23,$21
        x"02", x"B6", x"A8", x"20", -- ADD  $21,$21,$22
        x"32", x"D6", x"00", x"00", -- ANDI $22,$22,0 
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"D7", x"B0", x"25", -- OR   $22,$22,$23 
        x"AE", x"95", x"00", x"00", -- SW  $21,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        --10 
        x"32", x"F7", x"00", x"00", -- ANDI $23,$23,0
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"F5", x"B8", x"25", -- OR   $23,$23,$21
        x"02", x"B6", x"A8", x"20", -- ADD  $21,$21,$22
        x"32", x"D6", x"00", x"00", -- ANDI $22,$22,0 
        x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00",
        x"02", x"D7", x"B0", x"25", -- OR   $22,$22,$23
        x"AE", x"95", x"00", x"00", -- SW  $21,0($20)
        x"22", x"94", x"FF", x"FF", -- ADDI $20,$20,-1
        others => x"00");

begin
    process (addr) begin
        if (to_integer(unsigned(addr)) <= 1023) then
            d_out(31 downto 24) <= mem_array(to_integer(unsigned(addr)));
            if (to_integer(unsigned(addr))+1 <= 1023) then
                d_out(23 downto 16) <= mem_array(to_integer(unsigned(addr))+1);
                if (to_integer(unsigned(addr))+2 <= 1023) then
                    d_out(15 downto 8) <= mem_array(to_integer(unsigned(addr))+2);
                    if (to_integer(unsigned(addr))+3 <= 1023) then
                        d_out(7 downto 0) <= mem_array(to_integer(unsigned(addr))+3);
                    else d_out(7 downto 0) <= (others => '0'); end if;
                else d_out(15 downto 0) <= (others => '0'); end if;
            else d_out(23 downto 0) <= (others => '0'); end if;                    
        else d_out <= (others => '0');
        end if;
    end process;          
end;